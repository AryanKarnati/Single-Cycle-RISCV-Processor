module ControlUnit (
  input  logic [6:0] opcode,
  output logic       RegWrite,
  output logic       ALUSrc,
  output logic       MemWrite,
  output logic       MemToReg,
  output logic       Branch,
  output logic [1:0] ALUOp
);



always_comb begin
  // Default safe values
  RegWrite = 0;
  ALUSrc   = 0;
  MemWrite = 0;
  MemToReg = 0;
  Branch   = 0;
  ALUOp    = 2'b00;

  case (opcode)
    7'b0110011: begin // R-type
      RegWrite = 1;
      ALUSrc   = 0;
      MemToReg = 0;
      ALUOp    = 2'b10;
    end
    7'b0010011: begin // I-type (e.g., addi)
      RegWrite = 1;
      ALUSrc   = 1;
      MemToReg = 0;
      ALUOp    = 2'b00;
    end
    7'b0000011: begin // Load (e.g., lw)
      RegWrite = 1;
      ALUSrc   = 1;
      MemToReg = 1;
      ALUOp    = 2'b00;
    end
    7'b0100011: begin // Store (e.g., sw)
      RegWrite = 0;
      ALUSrc   = 1;
      MemWrite = 1;
      ALUOp    = 2'b00;
    end
    7'b1100011: begin // Branch (e.g., beq)
      RegWrite = 0;
      ALUSrc   = 0;
      Branch   = 1;
      ALUOp    = 2'b01;
    end
  endcase
end

endmodule

